//-----------------------------------------------------------------------------
// Copyright and license header
//
//-----------------------------------------------------------------------------
// File name: sif_driver_test.v
//-----------------------------------------------------------------------------
// Description:
//   TODO
//-----------------------------------------------------------------------------
// History:
//   - 2023-11-17 - federico g. zacchigna - Original version.
//
//-----------------------------------------------------------------------------




//-----------------------------------------------------------------------------
// Includes
//-----------------------------------------------------------------------------
//-----------------------------------------------------------------------------




//-----------------------------------------------------------------------------
// Module
//-----------------------------------------------------------------------------
module sif_driver_test #(
  // Word widths
  parameter I_WW = 6,
  parameter O_WW = 6
) (
  // clk, en, srst
  input             clk_i ,
  input             en_i  ,
  input             srst_i,
  // Input stream
  input  [I_WW-1:0] i_data_i,
  input             i_valid_i,
  output            i_ready_o,
  // Output stream
  output [O_WW-1:0] o_data_o,
  output            o_valid_o,
  input             o_ready_i
);
//-----------------------------------------------------------------------------
// Architecture
//-----------------------------------------------------------------------------

  //---------------------------------------------------------------------------
  // Constants
  //---------------------------------------------------------------------------
  localparam COUNTER_WIDTH = 16;
  localparam COUNTER_MAX   = 2**COUNTER_WIDTH-1;
  //---------------------------------------------------------------------------


  //---------------------------------------------------------------------------
  // Types
  //---------------------------------------------------------------------------
  //---------------------------------------------------------------------------


  //---------------------------------------------------------------------------
  // Signals
  //---------------------------------------------------------------------------
  // Control
  wire                     ien_s;
  reg  [COUNTER_WIDTH-1:0] counter_s;
  //---------------------------------------------------------------------------

  //---------------------------------------------------------------------------
  // Counter
  //---------------------------------------------------------------------------
  always @(posedge clk_i)
  begin
    if (srst_i) begin
      counter_s <= {COUNTER_WIDTH{1'b0}};
    end else if (ien_s) begin
      if (counter_s == COUNTER_MAX) begin
        counter_s <= {COUNTER_WIDTH{1'b0}};
      end else begin
        counter_s <= counter_s + {{COUNTER_WIDTH-1{1'b0}}, 1'b1};
      end
    end
  end
  //---------------------------------------------------------------------------


  //----------------------------------------------------------------------------
  // Stream Interface bypass
  //----------------------------------------------------------------------------
  assign ien_s     = 1'b1;
  assign o_data_o  = i_data_i;
  assign o_valid_o = i_valid_i;
  assign i_ready_o = o_ready_i;
  //----------------------------------------------------------------------------


  //----------------------------------------------------------------------------
  // Dump waves
  //----------------------------------------------------------------------------
  initial begin
    $dumpfile("waves.vcd");
    $dumpvars(1, sif_driver_test);
  end
  //----------------------------------------------------------------------------

endmodule
//------------------------------------------------------------------------------

